`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:49:26 05/17/2018 
// Design Name: 
// Module Name:    MatrixSumByMatrix 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MatrixSumByMatrix #(parameter N=100)(
	output [N-1:0]out);
	
assign out[12287:11904]=384'h0032fff200220036fff8002d002effee00060011006d0004fff8ff8fffe5000e002e0015ffc60045ffeffffd0006ffe5;
assign out[11903:11520]=384'hffe00056ffe2ffecffebffc6ffeb0001ffd2ff8f001d00220010004700020010ffc5ffd3000600290002ffc1ffec0023;
assign out[11519:11136]=384'hfff5fff60008ffa3fff8003affa1ffe0ffc6fffdfffffff4ffc6ffe20029ffffffda0006fff60046004e000b0013ffbe;
assign out[11135:10752]=384'hffc6fff8ffdb0009ffd0ffedffb6fff6ffdffff000510004000f0026002e0011fffcffaf000c0019ffc9ffefff9a0037;
assign out[10751:10368]=384'h000a0028ffdaffc3ffdc000e0009000b0059ffc5004efff4ffdafff8001b00420005000ffff7001b000c00050058ffaa;
assign out[10367:9984]=384'h0021fff8ffde005c000effc2ffdc002afffb007f002c0032ffd8000400280006ffd90032ffffffefffe8ffeaffe90028;
assign out[9983:9600]=384'hfff5ffc6ffd4003d003f00040036ffc6ffef002cffeb003bfff2ffac00040030ffd0ffbaffd6ffe1ffc5000a0017fff9;
assign out[9599:9216]=384'h004cffe30012ffca00100002001f0052ffd9003a00270060ffdc002e00210001003b0004001cffd9000bffdd002b0031;
assign out[9215:8832]=384'hffcf00090003ffcbff82002a000400000009ffe7ffc9ffd9ffcf003900000042000f001effbeffd10016ffd1ffee000a;
assign out[8831:8448]=384'hffc80013ffd3ffe30032fff6001a0002ffee001cffe3ffcc002bffb8ffdfffb00023ffe2006d0020ffc6ffe5ffdf000e;
assign out[8447:8064]=384'hfff5ffcafffcfff200160015fff9fff5ffa50022ffecffec002cfff9002cffb900020001ff7cffffffcc00430019000e;
assign out[8063:7680]=384'hffca0038001b003400010021ffc7ff7a000cfff50013fffbffef0001ffe0002e003effc7fffeffd1ffee0016ffd60024;
assign out[7679:7296]=384'hffdeffcfffdb000b00000059ffe900400015ffd50042ffd1000d0017ffaafffe002dffeb000b000bff9effd300060014;
assign out[7295:6912]=384'hffd1ffd700320000ffe1006e000d00090042002fffe20054ffd3fff70018002afff5fffbfffafff8ffbd001affc1ffde;
assign out[6911:6528]=384'h00010034000bffde000fffe40031ffcfffebffe4000e0002ffedffd0003cff8afff0ffe10004ffccffcc0009ff97fff8;
assign out[6527:6144]=384'hffd5ffcdffd5ffe1002e0032ffed003efffcffe8ffd3ffcaffb3ffbb0038fffa00230034fffeffc10018003affebffdb;
assign out[6143:5760]=384'hfff50006ffe9ffe6ffd10018000a0045001dffdc0061003b001b001a001d001e00060050004affe8fff700010029ffa7;
assign out[5759:5376]=384'hffe9001a0002ffe2fff9fff90000ffbeffef0009fffb004affb1ffffffacfffb0073ffd50025fff2ffc20024ffea0021;
assign out[5375:4992]=384'hffd6ff93001d0006ffe6fff3000effe0001400520022fffc002d0066003effd5000affef000c001500030032ffcc0001;
assign out[4991:4608]=384'h002a0020000fffe80006ffad0024002e0033003f000800380002fff0ffbc0004fff50032ffd40032002fffea0024ff9f;
assign out[4607:4224]=384'hffec000b0030ffe6fff6ffe6ffee0000003dffecffd0001dfff00036ffe2ffcaffdaffeeffea000e0080ffd9001d0060;
assign out[4223:3840]=384'h000affe8fff4ffe40041002cffe7002ffff2003f0088000d0026002a0017000efff8ffe8fff60007fff100170048ffb8;
assign out[3839:3456]=384'hffc00029ff9c005efff5001300030021ffd6ffe8000f00100000fffbffe0ffebffdc002700070007ffedffe5006affc5;
assign out[3455:3072]=384'hffe9ffc7ffd300010045ffe6ffc20044000effe8002a0007000cffbdffc6ffd70004fff4ffedffc800050035000b0067;
assign out[3071:2688]=384'hff8c00530003fff5ffffffd3003f0014001e00280015ffd2000500200022fff50002ffd9fff20007fffa005a0015ffbd;
assign out[2687:2304]=384'hfff3ffac0012ffc9ffd5fffc004100550003ffaaffebffec0008002dffecfffc0011ffc3ffc6ffedfffffff5000affaf;
assign out[2303:1920]=384'h0032001c001e0002ffe3000d0013ffdefff3fff5ffd1003fffd00074ffe7ffe5ffc1fffe001cffe5ffcc0034002bffb1;
assign out[1919:1536]=384'hffcb003800210001005200240036000c002a0009001a004c002bffe7001f00670005ffe4ffeeffab0009ffe800000006;
assign out[1535:1152]=384'hff9cffe900500025ffdc007b00120007ffdfffd4ffecffed0016002000190006002effce002d00100009fffffffc0022;
assign out[1151:768]=384'h002effd8ffb100360019001d004f000affe0ffcdffb10016fffdffc50001fff20022fff40009ffa1fffd001fffd1ffe3;
assign out[767:384]=384'hffdd001fffb80006ffd7ffccffd2ffc70001ffc1ffa7fff2ffebffe1ffb30020002d0004003a001bfffefffeffe2ffbc;
assign out[383:0]=384'hfff1000b001fffcfffed006e001dffd800410039fffe0043001300280047001e0007fff30049ffe2fff9ffc90021fffa;



endmodule
