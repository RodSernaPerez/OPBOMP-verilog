`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:07:33 05/17/2018 
// Design Name: 
// Module Name:    Pseudoinverses 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Pseudoinverses #(parameter N=100)(
	output [N-1:0]out);


assign out[38015:37632]=384'h0ff0f00f000fff0f00f000000ff0f00f000fff0f00f000000fa777053367780f286f25359bb5394610978a742fe8e414;
assign out[37631:37248]=384'h0000ff00f0000ff00fff0fff0000ff00f0000ff00fff0fef825cef4cf19422e44f5c2ee81bc30331b0b5c02d64e8afd1;
assign out[37247:36864]=384'h0f0f000ff0000fff0f00ff0f0f0f000ff0100fff0f00ef1f86f7e8d7d059606fab69f7877349f6a2c9ecce0e126613f6;
assign out[36863:36480]=384'hf0ff0f0fff00f0000f000000f1ff0f0fff00f0000f000000f01e1b7e5550d92229a3163058831bd81deab12dd8bca9ae;
assign out[36479:36096]=384'hf00fffffff00ff00fffffff0f00fffefff00ff00fffffef08c2eda9ffa93bd2b968dee9fca40c9e8f861c889dbe1b920;
assign out[36095:35712]=384'hff0fff00fff000fff0f00fffff0fff00fef001ffe0f00fffca6d8663e978e1a4c3be02baf8f6f4a021dcb5a75110052d;
assign out[35711:35328]=384'hff0f00fff0fff00ff0f00fffff0f00fff0fff00ff0f00fffc4498698f1eb9b4bb0966dfa1741fab11f0b8f7361c19409;
assign out[35327:34944]=384'h00fffffff000ff0000f00fff00fffffff000ff0000f00fff178bfdbe5436300259ebefb8c561da97724046f69ed97ed6;
assign out[34943:34560]=384'hf00ff0f0ffff0f00ff00f00ff00ff0f0ffff0f00ff00f00ff4521b02a7eb48534760f7bbd520d718fef8a0d9927c81a7;
assign out[34559:34176]=384'hf0f00fff0f000f00fff0fffff0e00fff0f000f00fff0ffff8161598d2f622d30aee6281d60c4c16398f67abc8ef7d8c0;
assign out[34175:33792]=384'hff00f0fff00f00f00ff0f0f0ff00f0fff00f00f00ff0f0f1ba3971a985efb7f96231fab0c9005b08565eb5868dd21eb6;
assign out[33791:33408]=384'hf00ffff0ff0ff00fff00fff0f01feff0ff0ff00ffe10ffe07215df29815e2af9df80c4d54c60b586079315e33dd1a07f;
assign out[33407:33024]=384'hf00fff000f00f00000f0000ff00fff000f00f00000f0001fe99bda305b2540417ca4902a795699d8f99a7e102c424a2a;
assign out[33023:32640]=384'h0fff00ffff0ff0f0ff00ff0f0ffe00ffff0ff0f0ff00ff0e6d9e3e6effe464ebf960996d3ff596a9a1ec0ac68b7a1623;
assign out[32639:32256]=384'hf0f0ff000f000f00fff0f00ff0e0ff001f000f00fff0f00ff4b32c859090c66a8ad3f81c31530a71ce16d91dbf997831;
assign out[32255:31872]=384'h0f00ff00f0f0ff0fff0f0f000f00ff00f1f0ff0fff0f0f00152b6b59e1a5dc6ccc0e79184a5d08365684352bd2d7036c;
assign out[31871:31488]=384'h00f000fff000ff00f000f0ff00f000fff000ff00f000f0ff3263443edf429e29e2a0114f4d5e91292f2c138bde0a0dc8;
assign out[31487:31104]=384'h00f00ff00000f00ff0ff0f0000f00ef00010f00ff1ff0f0057dcd9c44027e929730b1e43fc210ea17db992bf9fe36f90;
assign out[31103:30720]=384'h0f00ff0f00fffff0fffff0ff0f00ff0f00fffff0fffff0ff0935dc3a6e9ea06ed5adebd32b972799b584c96816ac26fe;
assign out[30719:30336]=384'hfff0000ffff0ff000f0fff00fff0000ffff1ff000f0fff0054a58a01d7e7b76205cb97818f16e42b7a31962ffc67acc5;
assign out[30335:29952]=384'h0ff00f00f00f0f0fffffff000ff01f00f00f0f0fffefff006e290be0472f5d6c1eac3e1ad96973cce122bb5bcbb6fa88;
assign out[29951:29568]=384'h000f000ff000f0f0000f0000000f000ff000f0f0000f0000532a71dc828c79492029909b83bfd69fa833c54ff517e8de;
assign out[29567:29184]=384'h0f0ff0f0f0000000000ff00f0e0ff0f1f0000010000ff00fdf1ba4a1816d418ccf5da69978da92cc1347b4a76395222e;
assign out[29183:28800]=384'h000f0ff000f0f00f0f0ffff0000f0ff101f0f00e0e0ffef0a01419e535d974518f3bc79a8dc54dfd1aa63f1f0a56398c;
assign out[28799:28416]=384'hfffff0ffff0ff000f0f0ff0ffffff0ffff0ff000f0f0ff0fbec8ba5fb71f9603f611ac1f21b89d49683057929c512f18;
assign out[28415:28032]=384'hf00ff00f00f0f0000fff0000f00fe00f00f0f0000fff0000dbc6107c92a1eb9898ccda3f6bfc6fb4abb955e34230ac62;
assign out[28031:27648]=384'hfff0ff0000fff0f0f00f0ffffff0ff0000eef0f0f00e0eff7a913cd422cf904dd83e56246ea6eb6c488da3d65769adff;
assign out[27647:27264]=384'hf00f0f0ff0000f0f0f0000f0f00f0f0ff0000f0f0f0000f08c086f5f9301b97c8f680483dd925638a6809a92e958b532;
assign out[27263:26880]=384'h0fff00000fffffffff00ff000fef00000ffffeffff10fe006cd807201abade6a8a8a7aadb436f6932111e45d436501c0;
assign out[26879:26496]=384'hfff00ff000ff0fff0f0ff0ffeff00ff000fe0fee0f0fe0ffa3fba3f13e6b0fb689b1c430f596c22a109409874417e504;
assign out[26495:26112]=384'h0ff0f0ffff0f000ffff0f0f00ff0f0ffff0f000ffff0f0f0ebe764b7390e5051df719ba62959446bd8e5f01eb157841e;
assign out[26111:25728]=384'hff0f000ff0f0f0ff0ff0f00fff0f100ff0f0f0ff1fe0f00f5d16461644abd0b50ec4a29cbfe0617636d0b148c3d474e2;
assign out[25727:25344]=384'hffffff00f0ff0f00f0fff000ffffff01f1fe0f00f0eff00033ebfb22a1cebdf303d8a77021a09719aeb0e5aafa8ccf63;
assign out[25343:24960]=384'hf0f000ff000ff0f00f0f0ffff0f000ff000ff0f00f0f0fff60d9818cf30c54f5fb1a2f9f3a1df1c8339bc5fed28fcf0b;
assign out[24959:24576]=384'h000f00ffff0f00f00f0fff00000f00ffff0f00f00e0fff001a9c46e3692a43682b3a4f58429ce0bf8810c9a919769ae0;
assign out[24575:24192]=384'hf000f0ffff000ffff0ff00f0f000e0feff000ffff0ff00f07729c360af3a25fddb8c3924fdbed98784ff75afe95bc541;
assign out[24191:23808]=384'h00ff00000f0ff0ffff0fffff00ef01000f0ff0ffff0fffff63bd20aa6bb5d38b9a6eaded07750850eacf997e516654f8;
assign out[23807:23424]=384'hff00f0ff0f0000f000ffffffff00f0ff0e0000f010ffefffeb60d46d6c95c8a323dd7d8d56781656473e5d0441f5e45b;
assign out[23423:23040]=384'hff0000f0f00ffff00ff0ff00ee0000f1f00fffe00ff0ff00bc4709307b03aad06beab3deb2fcb7b3f794129d3a53bf58;
assign out[23039:22656]=384'hff0ff00000f0ff00ff0000ffff0ff00000f0ff00ff0000ff5dbe898380b6bd41d78e35e4dc7d8d7697506833a4aeadee;
assign out[22655:22272]=384'h0fff00ff0000ff0ffffff0ff0fff00ff1000ff0ffffff0ff39ca1c2b35297ceccca220cfc06ecd9755b51c99b4ea816c;
assign out[22271:21888]=384'hff00f000f0f000f000fff0f0ff00f000f0f000f100fff0e08b77cc846a8c03213e7711e36f19fd927e450e8e06bfbb60;
assign out[21887:21504]=384'h00fff00fff00ff0fff00ffff00fff00fff00ff0fff00ffffe0ebe60bcc74dd80b5358ba7099f21f506b113056c2bb997;
assign out[21503:21120]=384'hf0ffff0f0f00ff0fff0f0ff0f0fffe0f0f00ff0fff0f0ff045eed87101506e098b004d466bb007beab4040b21f177dd0;
assign out[21119:20736]=384'hf00f0000f0ff0f0f00fff0f0f00f0000f0ff0f0f00fff0e07d8ac794dc2a82b1a8c41da3dddde55802b1ce02aea20bd7;
assign out[20735:20352]=384'hffff0ff0fffff0ff0fff000fffff0ff0fffff0ff0ffe000f63fdeffa9e887aad7ead741b6e86975d99f726a58ed98f52;
assign out[20351:19968]=384'hfffff0000fffff0f00f0f000fffff0000ffffe0f00f0f000608db3005eabc9e75692a84776febc1cc257c063cd1fd0e8;
assign out[19967:19584]=384'h00ff00f0ffffff00f00f00ff01ff01f0ffffff00f00f00ee80794199fae902bccefb67ed05e9d12fa9cf4eddc48a70d7;
assign out[19583:19200]=384'hf0fff00000f000f0f00f000ff0fff00000f010f0f00f000ff9a85a98a2e224a2d67e14b8bcd4b7521cba39fcdb12494b;
assign out[19199:18816]=384'hf0f0ff00ff000f0000fffffff0f0ff00ff200f0000fffffff184fc5193192f5e06cbfbda484649ff0c1a458394ba5e0f;
assign out[18815:18432]=384'hff0ffff00f00f00f000fff0fff0fffe00f00e00f001fff0ec37bcffd5c18e4c74f7ebe4cc23485fde259fb15b6917c6d;
assign out[18431:18048]=384'hf0fff0ff0000ffff0fff0000f0fff0ff0000ffff0fff000073fc65de30453e539cfa7702ff094570a667754200c55ee3;
assign out[18047:17664]=384'h0000000ffff0f0000f00fff00000000ffff0f0001f00fff04526b20fc66805361c944fe95b05c304ddb1160c75e0478b;
assign out[17663:17280]=384'hffffff0ff0000ff00f0ff0ffffffff0ef0000fe00f0fe0ffecf1d1497f3aabba8a2ea27c08d5874e724454e02224a4cd;
assign out[17279:16896]=384'hfff00fff000000f0000000f0fff00fff000000f0000000f0c5d56ddc62967de0133ca3c6e005a962f172a7debcb1cd6d;
assign out[16895:16512]=384'hff00f00ff000f00fff0ff0ffff00f00ff000f10fff0ff0ff93ec74a724439077e5172bfb614bb34b75c2bd3a538a8e55;
assign out[16511:16128]=384'hff0ffff000ff000f0ffff0ffff0efff001fe001f0ffff0efa30829e3ec8ee0553fcef0fae34ee102013ed41bf1e727b1;
assign out[16127:15744]=384'hf0ffff000000f000f0f0ff0ff0fffe000000f000f0f0ff0fd3b97d5a8851f550e770aa5a29b0701135eb154f5c16ac34;
assign out[15743:15360]=384'h000f000000f00ffff0ff0f0f000f000000f00ffff0ff0f0fcd698a2236ca9a5ea66e2f45a883967e32974a04f8db26e1;
assign out[15359:14976]=384'h0f000f0f00f0fff00f000fff0f000e0f00f0ffe00f011ffe433b4a3f34f638925fa8bfff03ce1df1f720c19ec0344fc4;
assign out[14975:14592]=384'hf0ff00fff000ffffffff0ff0f0ff00fff000ffffffff1ff0c5ef77acd00ffdf6d9cd5bf6d9de17f7180839f9af9b5f05;
assign out[14591:14208]=384'h0f0fff000fff000fffff0f000f0fff000fff000fffff0f012f2bd53569160578ff0d3c951aed6ebacca44b5fade005fb;
assign out[14207:13824]=384'hff0fffff0ff0f0f0f0000f00ff1fffff1ff0f1e0f0101f009b3a36bd6ff09482322e0a00bd7d384d88b9f138a93d0e34;
assign out[13823:13440]=384'hfff000f000000f00ffff000ffff000f000000f00ffff000fe9a1886c34931d1c42cd650b18ee231e4fc3d21d2fcfa226;
assign out[13439:13056]=384'h000ff0ff0000000ffff0ff0f000ff0ff0010000ffff0ef0f3224b0de047279e39c9cf6cc66c1e71e6a42eaecb9e3207a;
assign out[13055:12672]=384'h0fff0000f00f00f0000f000f0fff1000f00f00f0100f000e3dff35804dee3a606e873dfd33c5653f9252bb78320d5934;
assign out[12671:12288]=384'hfff00f00fff000fff00ff00ffff00f00fff000fff00ff00f1be418022ac406dca12571e93343fc91508214f3932e5f4e;
assign out[12287:11904]=384'hf0f00f000f0fff000ff0ff0ff1e00f000f0fff000ff0ff0fc47f7f78861bac193a55f864c71b2f2669aa3c45ea41381c;
assign out[11903:11520]=384'h00f0f0f0f0000ffff0000f0f00f1e1f0f0000ffff1000f0f1140d670abb5763146df89fd1f38f51d6f5c33533e6114ee;
assign out[11519:11136]=384'hffff0ff00f0fffff000f000fffff0ff00f0fffff000f000f67fb3b8517b7c7df0715145df2b6e7734969c3ea3804891c;
assign out[11135:10752]=384'h00f00ff0ffff0ffff0f0f0f000f00ff0ffff0ffff0f0f0f120ca7ca7ab9c2e958074adb086cb7f4e1becde030bd4c34b;
assign out[10751:10368]=384'h0fff00f000000ff00f0f0f000fff00f000010ff00e0f0f01283991c6ba645670ce267a2367f1dfa4bc0de60284b607b8;
assign out[10367:9984]=384'hf0f00fff000ff0f0fff0f00ff1f00fff000ff0f0fff0f00f918328eb59045a91f9b5f69fd79ed72803de8480108b02e8;
assign out[9983:9600]=384'hff0fff000f00f00f0f00f0ffef0fef000f00f00f0f00f0ffac1cdfa95e86e55a2854adbad5393a98d04b95551cea98df;
assign out[9599:9216]=384'hf00f0f00f0ff0f00f0ff00fff00f1f00f0ff1f00f0ff00fe6a9b0ac2d4d608e1f3a658feec009581a94c8553b3855c5e;
assign out[9215:8832]=384'hffff0f000ff00fff0ff00f0fffff0f000ff00fff0ff00f0fe38e1b244559adcd68c41e374165c13f0b48cad9df46da98;
assign out[8831:8448]=384'h0f0ff0000f0f00ff0fffff0f0f0ff0010f0f01ff0fffff0f0bb8ac311fea00b6b5177e4e75305284bd5600556e4f0cb3;
assign out[8447:8064]=384'hff0fff00fffff000ff0f0fffff0fff10fefef000ef0f0ffed96628268e8f132def0a7f8f0482d45099c2a399514955e8;
assign out[8063:7680]=384'h000f00000000f0fff00ff000000f00000000f0fff00ff0005586273113129dba41acd114029541bb1394a0de25b9d015;
assign out[7679:7296]=384'h00f0ff0ffff0f00f000ff0ff00f0ff0fffe0f00f000ff0ffb0b2833ad4f5744b2354efe33a53cd1e1741efc63a50e154;
assign out[7295:6912]=384'hf000f0fff00000f0fff0ff0ff000f0fff00000f0fff0ff0ed12da7d7d40c2f8398392ffc05e66fb2065f642a9f1a4ac0;
assign out[6911:6528]=384'hf00f0ff00f000ff0ff0ffff0f00f0ff00f000ff0ff0ffff063995feb59a3159cc85a9df2672ee286ab9734c615b098c4;
assign out[6527:6144]=384'hf0ff000f00f00000f0fffff0f0ff000f00f00000f0effff0eb88442bed6b903deaf3edf18f4efd3a6b33fa037b4aa711;
assign out[6143:5760]=384'hf000000fff0000000f0f0f0ff001101fff0000100f0f0f0fb27109387c5a35159446ed1deaf6b3fc1f6b1849561f2a5a;
assign out[5759:5376]=384'hf000f0f00f0000ff000f0ff0f000f0f00f0000ff000f0ff000560f581b35819371454aeadda224e67e306cebaf322543;
assign out[5375:4992]=384'hff000000ff0fff000f0000f0ef100000ef0eff100f0000f0ef07ed11dc66b81d1a8145e4697918bfdc489ac7eb181826;
assign out[4991:4608]=384'hff0ff00f0ff000000f00f00fff0ff11f0fe101000e01f00fa0ef3ad041314c08b47d623a541c2d2618730ac16bafd9f6;
assign out[4607:4224]=384'hfff0f00f0ff00ff0f00f00fffff0f00f0ff00ff0f00f00ff8e91fa9d16556eb1fa0914cc1c1bf94e9a4c44ac8f81466e;
assign out[4223:3840]=384'h00f00f0ff0f0f00f0ffff00000e00f0ff0f0f00f0ffef000a2e8494f72898188127e87604818587ade47ea41c3219f12;
assign out[3839:3456]=384'h0f000000fffffff00f0f0fff1e000000fffffef00f0f0fef3f274097a9c3cae1b8dc5aca7cbfcc5f71ea6823fd186dd0;
assign out[3455:3072]=384'hfff0f0fffff0f0f00f000ffffff0f0ffffe0f0f00f000fffbcc564ddcbd6519a265768dff94f73a55f79e10cff66752b;
assign out[3071:2688]=384'h00ffffff0fff0fff00f000ff00fffeff0fff0eff10f000ff06a85ab266e92c79118a8af5c658a7c9e46589074c60995d;
assign out[2687:2304]=384'hf0f00fffffff00f0f00ffffff0e00fffffff00f0f12feffe3f72c919e374690593104f59c554ae3921921c57319804b4;
assign out[2303:1920]=384'hfffff00f00f000f0ffff0ffffffff00e00f000f0ffff0fffa7b4d94dc4d947e2e9df4bf817bbf4b0f3e7901b252dbfca;
assign out[1919:1536]=384'hf00ff0000000f000000ffff0f00ff0000000f010000ffff0e7d5b445612b53053870a789102775c323b6ebeff069da97;
assign out[1535:1152]=384'h000000f0f0ff00000f00ff0f000001f0f0ff00000f10ff1f582a19e5ffeee1a00a88ca7c37381fd57ffe523ca5e2d4b8;
assign out[1151:768]=384'h0f0ffff00f00fffffff0f0f00f0ffff00f00fffffff0f0f0193d3e41fd844eaaec4b45c16bf43cef9b882974f99dec9e;
assign out[767:384]=384'hf00ffff0f0ff0ff0f00ffff0f00fffe0f0ff0ff0f00ffff04375acd269beb839513a4bc32241f0245b2d789d95ba361b;
assign out[383:0]=384'h0f000f000ff00ffff0ff0fff0e000f010ff01ffff0ff0fffa852674275d937ea6a4627598d1160db110bd1f2a4625cdf;

endmodule
